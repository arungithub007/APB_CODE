class apb_seq_item extends uvm_sequence_item;// transaction
  
  //we have to declare data signals and control fields
  rand bit        	    [7:0] paddr;
  rand bit                    pwrite;
       bit                    psel;
       bit                    penable;
  rand bit        	   [31:0] pwdata;
       bit        	   [31:0] prdata;
       bit                    pready;
  
  `uvm_object_utils_begin(apb_seq_item)
  `uvm_field_int(paddr,UVM_ALL_ON)
  `uvm_field_int(pwrite,UVM_ALL_ON)
  `uvm_field_int(psel,UVM_ALL_ON)
  `uvm_field_int(penable,UVM_ALL_ON)
  `uvm_field_int(pwdata,UVM_ALL_ON)
  `uvm_field_int(prdata,UVM_ALL_ON) 
  `uvm_field_int(pready,UVM_ALL_ON) 
  `uvm_object_utils_end


  //constructor new
  function new(string name="apb_seq_item");
    super.new(name);
  endfunction:new
  
 endclass:apb_seq_item
